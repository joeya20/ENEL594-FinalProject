module simple3;

logic test;

endmodule